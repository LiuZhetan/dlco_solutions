module Hex2Segcode (
    input [3:0] x,
    output [7:0] y
);
    wire [3:0] key;
    wire [7:0] out;
    assign key = x;
    assign y = out;
    MuxKeyWithDefault #(16, 4, 8) mutex (out, key, 8'b1, {
    4'h0, ~(8'b11111100),
    4'h1, ~(8'b01100000),
    4'h2, ~(8'b11011010),
    4'h3, ~(8'b11110010),
    4'h4, ~(8'b01100110),
    4'h5, ~(8'b10110110),
    4'h6, ~(8'b10111110),
    4'h7, ~(8'b11100000),
    4'h8, ~(8'b11111110),
    4'h9, ~(8'b11100110),
    4'ha, ~(8'b11101110),
    4'hb, ~(8'b00111110),
    4'hc, ~(8'b00011010),
    4'hd, ~(8'b01111010),
    4'he, ~(8'b11011110),
    4'hf, ~(8'b10001110)
  });
endmodule